library ieee;
use IEEE.std_logic_1164.all;

entity fulladder is
    port(
        fa_in0         : in std_logic;
        fa_in1         : in std_logic;
        fa_carry_in    : in std_logic;
        fa_carry_out   : out std_logic;
        fa_output      : out std_logic
    );
end fulladder;

architecture structural of fulladder is
    --Declare component for structural modeling
    component halfadder is
        port(
           a            : in std_logic;
           b            : in std_logic;
           c            : out std_logic;
           sum          : out std_logic             
        );
    end component;
    
    component orgate is
        port(
            x           : in std_logic;
            y           : in std_logic;
            z           : out std_logic       
        );
    end component;
    
    --Initialize signal
    signal sum0         : std_logic;
    signal sum1         : std_logic;
    signal sum2         : std_logic;
    
    --Connecting components to make a 2 bit full adder
    begin
        u1      :   halfadder port map (a => fa_in0, b => fa_in1, c => sum1, sum => sum0);
        u2      :   halfadder port map (a => sum0,b => fa_carry_in, c => sum2, sum => fa_output);
        u3      :   orgate    port map (x => sum2, y => sum1, z => fa_carry_out);
end structural;
