library IEEE;
use IEEE.STD_LOGIC_1164.ALL; -- STD_LOGIC and STD_LOGIC_VECTOR
use IEEE.numeric_std.ALL; -- to_integer and unsigned

entity registers is
-- This component is described in the textbook, starting on section 4.3 
-- The indices of each of the registers can be found on the LEGv8 Green Card
-- Keep in mind that register 31 (XZR) has a constant value of 0 and cannot be overwritten
-- This should only write on the negative edge of Clock when RegWrite is asserted.
-- Reads should be purely combinatorial, i.e. they don't depend on Clock
-- HINT: Use the provided dmem.vhd as a starting point
port(RR1      : in  STD_LOGIC_VECTOR (4 downto 0); 
     RR2      : in  STD_LOGIC_VECTOR (4 downto 0); 
     WR       : in  STD_LOGIC_VECTOR (4 downto 0); 
     WD       : in  STD_LOGIC_VECTOR (63 downto 0);
     RegWrite : in  STD_LOGIC;
     Clock    : in  STD_LOGIC;
     RD1      : out STD_LOGIC_VECTOR (63 downto 0);
     RD2      : out STD_LOGIC_VECTOR (63 downto 0);
     --Probe ports used for testing.
     -- Notice the width of the port means that you are 
     --      reading only part of the register file. 
     -- This is only for debugging
     -- You are debugging a sebset of registers here
     -- Temp registers: $X9 & $X10 & X11 & X12 
     -- 4 refers to number of registers you are debugging
     DEBUG_TMP_REGS : out STD_LOGIC_VECTOR(64*4 - 1 downto 0);
     -- Saved Registers X19 & $X20 & X21 & X22 
     DEBUG_SAVED_REGS : out STD_LOGIC_VECTOR(64*4 - 1 downto 0)
);
end registers;

architecture behavioral of registers is
     type ByteArray is array(0 to 32) of STD_LOGIC_VECTOR(63 downto 0);
     signal reg: ByteArray;
begin
     process(Clock, RR1, RR2, WR, WD, RegWrite)
          variable addrW:integer;
          variable addrR1:integer;
          variable addrR2: integer;
          variable first:boolean := true; --Initialization
     begin
          if(first) then           --Initilize the value of the register
               --Temp Register
               reg(9)  <= X"0000000000000000";
               reg(10) <= X"0000000000000001";
               reg(11) <= X"0000000000000002";
               reg(12) <= X"0000000000000004";
               reg(13) <= X"0000000000000008";
               reg(14) <= X"0000000000000010";
               reg(15) <= X"0000000000000020";

               --Saved register
               reg(19) <= X"0000000000000008";
               reg(20) <= X"0000000000000000";
               reg(21) <= X"0000000000000002";
               reg(22) <= X"0000000000000004";
               reg(23) <= X"0000000000000010";
               reg(24) <= X"0000000000000020";
               reg(25) <= X"0000000000000040";
               reg(26) <= X"0000000000000080";
               reg(27) <= X"0000000000000080";
               
               first := false;
          end if;
          
          --Write process
          if Clock = '0' and Clock'event and RegWrite='1' then
               addrW := to_integer(unsigned(WR));
               reg(addrW) <= WD;
               if addrW = 0 or addrW = 31 then report "XZR cannot be overwrite"
                    severity error;
               end if;
          end if;

          --Read process          
          addrR1 := to_integer(unsigned(RR1));
          addrR2 := to_integer(unsigned(RR2));

          RD1 <= reg(addrR1);
          RD2 <= reg(addrR2);
     end process;

end behavioral;
