library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_imem is
    --Declare entity
end tb_imem;

architecture behavioral of tb_imem is
    component imem is
        port(
            Address  : in  STD_LOGIC_VECTOR(63 downto 0); -- Address to read from
            ReadData : out STD_LOGIC_VECTOR(31 downto 0)
        );
    end component;

    signal tb_Address : STD_LOGIC_VECTOR(63 downto 0);
    signal tb_ReadData: STD_LOGIC_VECTOR(31 downto 0);

begin
    uut: imem port map(Address => tb_Address, ReadData => tb_ReadData);

    stimulus: process
    begin
        tb_Address <= (others=>'0');
        wait for 500 ns;
    end process;
end behavioral;
